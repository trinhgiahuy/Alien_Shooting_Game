--* ><(((('> * Puli puli * ><(((('> // Ƹ̵̡Ӝ̵̨̄Ʒ * swish swish* Ƹ̵̡Ӝ̵̨̄Ʒ Ƹ̵̡Ӝ̵̨̄Ʒ // (っ◕‿◕)╭∩╮^H^H^Hっ
LIBRARY ieee;USE ieee.std_logic_1164.all;USE ieee.std_logic_arith.all;ENTITY z_black_box IS PORT(clk:IN std_logic;color_BGR:IN std_logic_vector(23 DOWNTO 0);rst_n:IN std_logic;x_coord:IN std_logic_vector(7 DOWNTO 0);y_coord:IN std_logic_vector(7 DOWNTO 0);if_you_name:OUT std_logic_vector(7 DOWNTO 0);iotre_will:OUT std_logic;like_this:OUT std_logic;of_this_course:OUT std_logic;throw_you_out:OUT std_logic;your_signals:OUT std_logic);END z_black_box ;LIBRARY ieee;USE ieee.std_logic_1164.all;USE ieee.std_logic_arith.all;LIBRARY pre_made;ARCHITECTURE struct OF z_black_box IS SIGNAL zf54907441:std_logic;SIGNAL frame_done:std_logic;SIGNAL z3417d2827:std_logic_vector(23 DOWNTO 0);SIGNAL write:std_logic;SIGNAL z187d0b354:std_logic_vector(7 DOWNTO 0);SIGNAL z88ece3df0:std_logic_vector(7 DOWNTO 0);COMPONENT z_black_box_p PORT(z9544d0e66:IN std_logic_vector(7 DOWNTO 0);zf54907441:IN std_logic ;z5efa2601c:IN std_logic_vector(7 DOWNTO 0);zd1385ccb0:IN std_logic_vector(23 DOWNTO 0);clk:IN std_logic ;rst_n:IN std_logic ;frame_done:OUT std_logic ;z3417d2827:OUT std_logic_vector(23 DOWNTO 0);write:OUT std_logic ;z187d0b354:OUT std_logic_vector(7 DOWNTO 0);z88ece3df0:OUT std_logic_vector(7 DOWNTO 0));END COMPONENT;COMPONENT z_black_box_y PORT(clk:IN std_logic ;color_BGR:IN std_logic_vector(23 DOWNTO 0);frame_done:IN std_logic ;rst_n:IN std_logic ;write:IN std_logic ;x_coord:IN std_logic_vector(7 DOWNTO 0);y_coord:IN std_logic_vector(7 DOWNTO 0);if_you_name:OUT std_logic_vector(7 DOWNTO 0);iotre_will:OUT std_logic ;like_this:OUT std_logic ;of_this_course:OUT std_logic ;throw_you_out:OUT std_logic ;w_rdy:OUT std_logic ;your_signals:OUT std_logic);END COMPONENT;FOR ALL:z_black_box_p USE ENTITY pre_made.z_black_box_p;FOR ALL:z_black_box_y USE ENTITY pre_made.z_black_box_y;BEGIN U_1:z_black_box_p PORT MAP(z9544d0e66=>x_coord,zf54907441=>zf54907441,z5efa2601c=>y_coord,zd1385ccb0=>color_BGR,clk=>clk,rst_n=>rst_n,frame_done=>frame_done,z3417d2827=>z3417d2827,write=>write,z187d0b354=>z187d0b354,z88ece3df0=>z88ece3df0);U_0:z_black_box_y PORT MAP(clk=>clk,color_BGR=>z3417d2827,frame_done=>frame_done,rst_n=>rst_n,write=>write,x_coord=>z187d0b354,y_coord=>z88ece3df0,if_you_name=>if_you_name,iotre_will=>iotre_will,like_this=>like_this,of_this_course=>of_this_course,throw_you_out=>throw_you_out,w_rdy=>zf54907441,your_signals=>your_signals);END struct;