--* ><(((('> * Puli puli * ><(((('> // Ƹ̵̡Ӝ̵̨̄Ʒ * swish swish* Ƹ̵̡Ӝ̵̨̄Ʒ Ƹ̵̡Ӝ̵̨̄Ʒ // (っ◕‿◕)╭∩╮^H^H^Hっ
LIBRARY ieee;USE ieee.std_logic_1164.all;USE ieee.std_logic_arith.all;ENTITY z_black_box_s IS PORT(clk:IN std_logic;rst_n:IN std_logic;z7f53ee971:IN std_logic;zea9c5ae7c:OUT std_logic;z7975aa26e:OUT std_logic;z2ebb22097:OUT std_logic);END z_black_box_s ;LIBRARY ieee;USE ieee.std_logic_1164.all;USE ieee.std_logic_arith.all;ARCHITECTURE fsm OF z_black_box_s IS SIGNAL z009e7c1f9:std_logic_vector(17 DOWNTO 0);SIGNAL zedc5ef274:integer RANGE 10 DOWNTO 0;SIGNAL zbddb18e97:integer RANGE 17 DOWNTO 0;TYPE STATE_TYPE IS(z300f5740b,z82451b49a,z5b4a4026f,z3d9d4ca12,z57e441642,ze7b757c44);SIGNAL zdf0be1ce6:STATE_TYPE;SIGNAL ze8e79043b:STATE_TYPE;BEGIN z9149816e0:PROCESS(clk,rst_n)BEGIN IF(rst_n='0')THEN zdf0be1ce6<=z300f5740b;z009e7c1f9<="111011111111001110";zedc5ef274<=0;zbddb18e97<=17;ELSIF(clk'EVENT AND clk='1')THEN zdf0be1ce6<=ze8e79043b;CASE zdf0be1ce6 IS WHEN z5b4a4026f=>zbddb18e97<=zbddb18e97-1;WHEN ze7b757c44=>zedc5ef274<=zedc5ef274 + 1;zbddb18e97<=17;WHEN OTHERS=>NULL;END CASE;END IF;END PROCESS z9149816e0;z145fbcc0d:PROCESS(zedc5ef274,zdf0be1ce6,zbddb18e97,z7f53ee971)BEGIN CASE zdf0be1ce6 IS WHEN z300f5740b=>IF(z7f53ee971='1')THEN ze8e79043b<=z82451b49a;ELSE ze8e79043b<=z300f5740b;END IF;WHEN z82451b49a=>IF(z7f53ee971='0')THEN ze8e79043b<=z3d9d4ca12;ELSE ze8e79043b<=z82451b49a;END IF;WHEN z5b4a4026f=>ze8e79043b<=z300f5740b;WHEN z3d9d4ca12=>IF(z7f53ee971='1'AND zbddb18e97=0)THEN ze8e79043b<=ze7b757c44;ELSIF(z7f53ee971='1')THEN ze8e79043b<=z5b4a4026f;ELSE ze8e79043b<=z3d9d4ca12;END IF;WHEN z57e441642=>ze8e79043b<=z57e441642;WHEN ze7b757c44=>IF(zedc5ef274=7)THEN ze8e79043b<=z57e441642;ELSE ze8e79043b<=z300f5740b;END IF;WHEN OTHERS=>ze8e79043b<=z300f5740b;END CASE;END PROCESS z145fbcc0d;z822bdb2c3:PROCESS(z009e7c1f9,zdf0be1ce6,zbddb18e97)BEGIN zea9c5ae7c<='0';z7975aa26e<='0';z2ebb22097<='0';CASE zdf0be1ce6 IS WHEN z300f5740b=>zea9c5ae7c<=z009e7c1f9(zbddb18e97);WHEN z82451b49a=>zea9c5ae7c<=z009e7c1f9(zbddb18e97);z2ebb22097<='1';WHEN z3d9d4ca12=>zea9c5ae7c<=z009e7c1f9(zbddb18e97);WHEN z57e441642=>z7975aa26e<='1';WHEN OTHERS=>NULL;END CASE;END PROCESS z822bdb2c3;END fsm;