--* ><(((('> * Puli puli * ><(((('> // Ƹ̵̡Ӝ̵̨̄Ʒ * swish swish* Ƹ̵̡Ӝ̵̨̄Ʒ Ƹ̵̡Ӝ̵̨̄Ʒ // (っ◕‿◕)╭∩╮^H^H^Hっ
LIBRARY ieee;USE ieee.std_logic_1164.all;USE ieee.std_logic_arith.all;ENTITY z_black_box_k IS PORT(clk:IN std_logic;zf1caf1a47:IN std_logic_vector(23 DOWNTO 0);rst_n:IN std_logic;z28f400601:IN std_logic;write:IN std_logic;zdf77ec582:IN std_logic_vector(7 DOWNTO 0);z187d0b354:IN std_logic_vector(7 DOWNTO 0);z5e19774c6:IN std_logic_vector(7 DOWNTO 0);z88ece3df0:IN std_logic_vector(7 DOWNTO 0);z3417d2827:OUT std_logic_vector(23 DOWNTO 0);w_rdy:OUT std_logic);END z_black_box_k ;LIBRARY ieee;USE ieee.std_logic_1164.all;USE ieee.std_logic_arith.all;LIBRARY pre_made;ARCHITECTURE struct OF z_black_box_k IS SIGNAL z98552069b:std_logic;SIGNAL ze72d2c2a4:std_logic_vector(7 DOWNTO 0);SIGNAL z508ec0017:std_logic;SIGNAL zb48298c48:std_logic;SIGNAL z9f041aaff:std_logic;SIGNAL zcf058ee7c:std_logic;SIGNAL z75dc1577a:std_logic_vector(7 DOWNTO 0);SIGNAL z833ab3bd5:std_logic_vector(7 DOWNTO 0);SIGNAL zc57c46db4:std_logic_vector(7 DOWNTO 0);SIGNAL z1ea89dc0d:std_logic_vector(7 DOWNTO 0);SIGNAL zcd48e1f4f:std_logic_vector(7 DOWNTO 0);SIGNAL z36424fa31:std_logic_vector(7 DOWNTO 0);SIGNAL z0068e7d64:std_logic_vector(7 DOWNTO 0);SIGNAL zb30429bb4:std_logic_vector(7 DOWNTO 0);SIGNAL z28c1a03db:std_logic;SIGNAL z921c03197:std_logic_vector(23 DOWNTO 0);SIGNAL zb488040b4:std_logic_vector(23 DOWNTO 0);SIGNAL z2677755d9:std_logic_vector(7 DOWNTO 0);SIGNAL z00b23bf66:std_logic_vector(7 DOWNTO 0);SIGNAL zaaac8007d:std_logic_vector(7 DOWNTO 0);SIGNAL zd4810c102:std_logic_vector(7 DOWNTO 0);COMPONENT z_black_box_f PORT(clk:IN std_logic ;zceb2b781a:IN std_logic ;rst_n:IN std_logic ;z98552069b:OUT std_logic ;z28c1a03db:OUT std_logic ;w_rdy:OUT std_logic);END COMPONENT;COMPONENT z_black_box_w PORT(clk:IN std_logic ;z28c1a03db:IN std_logic ;zd58ce0c39:IN std_logic_vector(23 DOWNTO 0);rst_n:IN std_logic ;write:IN std_logic ;z2677755d9:IN std_logic_vector(7 DOWNTO 0);zaaac8007d:IN std_logic_vector(7 DOWNTO 0);z921c03197:OUT std_logic_vector(23 DOWNTO 0));END COMPONENT;FOR ALL:z_black_box_f USE ENTITY pre_made.z_black_box_f;FOR ALL:z_black_box_w USE ENTITY pre_made.z_black_box_w;BEGIN z508ec0017<=z28c1a03db AND z98552069b;zb48298c48<=z28c1a03db AND NOT(z98552069b);z75dc1577a<=z187d0b354 AND ze72d2c2a4;z833ab3bd5<=NOT(ze72d2c2a4)AND zdf77ec582;zc57c46db4<=z88ece3df0 AND ze72d2c2a4;z1ea89dc0d<=NOT(ze72d2c2a4)AND z5e19774c6;zcd48e1f4f<=z187d0b354 AND NOT(ze72d2c2a4);z36424fa31<=ze72d2c2a4 AND zdf77ec582;z0068e7d64<=z88ece3df0 AND NOT(ze72d2c2a4);zb30429bb4<=ze72d2c2a4 AND z5e19774c6;z9f041aaff<=NOT(z98552069b)AND write;zcf058ee7c<=write AND z98552069b;ze72d2c2a4<=z98552069b & z98552069b & z98552069b & z98552069b & z98552069b & z98552069b & z98552069b & z98552069b;z33254a172:PROCESS(z921c03197, zb488040b4, z98552069b)BEGIN CASE z98552069b IS WHEN'0'=>z3417d2827<=z921c03197;WHEN'1'=>z3417d2827<=zb488040b4;WHEN OTHERS=>z3417d2827<=(OTHERS=>'X');END CASE;END PROCESS z33254a172;z2677755d9<=z75dc1577a OR z833ab3bd5;z00b23bf66<=zcd48e1f4f OR z36424fa31;zaaac8007d<=zc57c46db4 OR z1ea89dc0d;zd4810c102<=z0068e7d64 OR zb30429bb4;U_2:z_black_box_f PORT MAP(clk=>clk,zceb2b781a=>z28f400601,rst_n=>rst_n,z98552069b=>z98552069b,z28c1a03db=>z28c1a03db,w_rdy=>w_rdy);U_0:z_black_box_w PORT MAP(clk=>clk,z28c1a03db=>z508ec0017,zd58ce0c39=>zf1caf1a47,rst_n=>rst_n,write=>zcf058ee7c,z2677755d9=>z2677755d9,zaaac8007d=>zaaac8007d,z921c03197=>z921c03197);U_1:z_black_box_w PORT MAP(clk=>clk,z28c1a03db=>zb48298c48,zd58ce0c39=>zf1caf1a47,rst_n=>rst_n,write=>z9f041aaff,z2677755d9=>z00b23bf66,zaaac8007d=>zd4810c102,z921c03197=>zb488040b4);END struct;