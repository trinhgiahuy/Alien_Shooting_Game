--* ><(((('> * Puli puli * ><(((('> // Ƹ̵̡Ӝ̵̨̄Ʒ * swish swish* Ƹ̵̡Ӝ̵̨̄Ʒ Ƹ̵̡Ӝ̵̨̄Ʒ // (っ◕‿◕)╭∩╮^H^H^Hっ
LIBRARY ieee;USE ieee.std_logic_1164.all;USE ieee.std_logic_arith.all;ENTITY mem_ctl_block IS PORT(clk:IN std_logic;pixd_w_done:IN std_logic;rst_n:IN std_logic;banksel:OUT std_logic;nullify:OUT std_logic;w_rdy:OUT std_logic);END mem_ctl_block ;LIBRARY ieee;USE ieee.std_logic_1164.all;USE ieee.std_logic_arith.all;ARCHITECTURE fsm OF mem_ctl_block IS TYPE STATE_TYPE IS(z77ca48e55,zd561de642,zfbdccd934,z0f0974e71);SIGNAL zdf0be1ce6:STATE_TYPE;SIGNAL ze8e79043b:STATE_TYPE;SIGNAL ze03a9bfed:std_logic ;SIGNAL z0650cbe3e:std_logic ;BEGIN z9149816e0:PROCESS(clk,rst_n)BEGIN IF(rst_n='0')THEN zdf0be1ce6<=z77ca48e55;ze03a9bfed<='0';z0650cbe3e<='0';ELSIF(clk'EVENT AND clk='1')THEN zdf0be1ce6<=ze8e79043b;CASE zdf0be1ce6 IS WHEN zd561de642=>ze03a9bfed<=not ze03a9bfed;WHEN zfbdccd934=>z0650cbe3e<='1';WHEN z0f0974e71=>z0650cbe3e<='0';WHEN OTHERS=>NULL;END CASE;END IF;END PROCESS z9149816e0;z145fbcc0d:PROCESS(zdf0be1ce6,pixd_w_done)BEGIN CASE zdf0be1ce6 IS WHEN z77ca48e55=>IF(pixd_w_done='1')THEN ze8e79043b<=zd561de642;ELSE ze8e79043b<=z77ca48e55;END IF;WHEN zd561de642=>ze8e79043b<=zfbdccd934;WHEN zfbdccd934=>ze8e79043b<=z0f0974e71;WHEN z0f0974e71=>IF(pixd_w_done='0')THEN ze8e79043b<=z77ca48e55;ELSE ze8e79043b<=z0f0974e71;END IF;WHEN OTHERS=>ze8e79043b<=z77ca48e55;END CASE;END PROCESS z145fbcc0d;z822bdb2c3:PROCESS(zdf0be1ce6)BEGIN w_rdy<='0';CASE zdf0be1ce6 IS WHEN z77ca48e55=>w_rdy<='1';WHEN OTHERS=>NULL;END CASE;END PROCESS z822bdb2c3;banksel<=ze03a9bfed;nullify<=z0650cbe3e;END fsm;