--* ><(((('> * Puli puli * ><(((('> // Ƹ̵̡Ӝ̵̨̄Ʒ * swish swish* Ƹ̵̡Ӝ̵̨̄Ʒ Ƹ̵̡Ӝ̵̨̄Ʒ // (っ◕‿◕)╭∩╮^H^H^Hっ
LIBRARY ieee;USE ieee.std_logic_1164.all;USE ieee.std_logic_arith.all;ENTITY debounce IS PORT(btn:IN std_logic_vector(3 DOWNTO 0);clk:IN std_logic;rst_n:IN std_logic;deb_btn:OUT std_logic_vector(3 DOWNTO 0));END debounce ;LIBRARY ieee;USE ieee.std_logic_1164.all;USE ieee.std_logic_arith.all;ARCHITECTURE struct OF debounce IS SIGNAL z0068e7d64:std_logic_vector(3 DOWNTO 0);SIGNAL z269042a3a:std_logic_vector(3 DOWNTO 0);SIGNAL z4fd12da22:std_logic_vector(3 DOWNTO 0);SIGNAL zc82b72865:std_logic_vector(3 DOWNTO 0);SIGNAL zce55af2db:std_logic_vector(3 DOWNTO 0);SIGNAL z2ed06566a:std_logic_vector(3 DOWNTO 0);SIGNAL zaa248e088:std_logic_vector(3 DOWNTO 0);SIGNAL zd144acfdd:std_logic_vector(3 DOWNTO 0);SIGNAL z48d1fd67d:std_logic_vector(3 DOWNTO 0);SIGNAL z65c50f750:std_logic_vector(3 DOWNTO 0);SIGNAL z99d1d6516:std_logic_vector(3 DOWNTO 0);SIGNAL zde1de9e8b:std_logic_vector(3 DOWNTO 0);SIGNAL z13563f2fa:std_logic_vector(3 DOWNTO 0);BEGIN z269042a3a<=z48d1fd67d;zce55af2db<=NOT(z48d1fd67d);zba7bd6dd5:PROCESS(clk, rst_n)BEGIN IF(rst_n='0')THEN z48d1fd67d<="0000";ELSIF(clk'EVENT AND clk='1')THEN z48d1fd67d<=z0068e7d64;END IF;END PROCESS zba7bd6dd5;z4fd12da22<=z65c50f750;z2ed06566a<=NOT(z65c50f750);zc9774e8a0:PROCESS(clk, rst_n)BEGIN IF(rst_n='0')THEN z65c50f750<="0000";ELSIF(clk'EVENT AND clk='1')THEN z65c50f750<=z269042a3a;END IF;END PROCESS zc9774e8a0;zc82b72865<=z99d1d6516;zaa248e088<=NOT(z99d1d6516);zd61aa8882:PROCESS(clk, rst_n)BEGIN IF(rst_n='0')THEN z99d1d6516<="0000";ELSIF(clk'EVENT AND clk='1')THEN z99d1d6516<=z4fd12da22;END IF;END PROCESS zd61aa8882;zd144acfdd<=NOT(zde1de9e8b);z71eb9a290:PROCESS(clk, rst_n)BEGIN IF(rst_n='0')THEN zde1de9e8b<="0000";ELSIF(clk'EVENT AND clk='1')THEN zde1de9e8b<=btn;END IF;END PROCESS z71eb9a290;deb_btn<=z13563f2fa;z61d5e22f5:PROCESS(clk, rst_n)BEGIN IF(rst_n='0')THEN z13563f2fa<="0000";ELSIF(clk'EVENT AND clk='1')THEN z13563f2fa<=zc82b72865;END IF;END PROCESS z61d5e22f5;z0068e7d64<=btn AND zaa248e088 AND z2ed06566a AND zce55af2db AND zd144acfdd;END struct;