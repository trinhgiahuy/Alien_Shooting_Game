--* ><(((('> * Puli puli * ><(((('> // Ƹ̵̡Ӝ̵̨̄Ʒ * swish swish* Ƹ̵̡Ӝ̵̨̄Ʒ Ƹ̵̡Ӝ̵̨̄Ʒ // (っ◕‿◕)╭∩╮^H^H^Hっ
LIBRARY ieee;USE ieee.std_logic_1164.all;USE ieee.std_logic_arith.all;ENTITY z_black_box_w IS PORT(clk:IN std_logic;z28c1a03db:IN std_logic;zd58ce0c39:IN std_logic_vector(23 DOWNTO 0);rst_n:IN std_logic;write:IN std_logic;z2677755d9:IN std_logic_vector(7 DOWNTO 0);zaaac8007d:IN std_logic_vector(7 DOWNTO 0);z921c03197:OUT std_logic_vector(23 DOWNTO 0));END z_black_box_w ;LIBRARY ieee;USE ieee.std_logic_1164.all;USE ieee.std_logic_arith.all;LIBRARY pre_made;ARCHITECTURE struct OF z_black_box_w IS SIGNAL z508ec0017:std_logic;SIGNAL z1934d98a3:std_logic;SIGNAL zb48298c48:std_logic;SIGNAL z9f041aaff:std_logic;SIGNAL zcf058ee7c:std_logic;SIGNAL ze6d31b4ac:std_logic;SIGNAL z1b791bfd5:std_logic;SIGNAL z45a1dff88:std_logic;SIGNAL zc83e54d35:std_logic_vector(2 DOWNTO 0);SIGNAL z22f92b4dd:std_logic;SIGNAL z75dc1577a:std_logic;SIGNAL z833ab3bd5:std_logic;SIGNAL zc57c46db4:std_logic;SIGNAL z1ea89dc0d:std_logic;SIGNAL zcd48e1f4f:std_logic;SIGNAL z36424fa31:std_logic;SIGNAL z0068e7d64:std_logic;SIGNAL zb30429bb4:std_logic;SIGNAL z36f79a239:std_logic_vector(3 DOWNTO 0);SIGNAL z3417d2827:std_logic_vector(23 DOWNTO 0);SIGNAL z564ee05a3:std_logic_vector(23 DOWNTO 0);SIGNAL z0a9315da3:std_logic_vector(23 DOWNTO 0);SIGNAL z6bb6c7052:std_logic_vector(23 DOWNTO 0);SIGNAL z163c5325c:std_logic_vector(23 DOWNTO 0);SIGNAL z84b2eb77e:std_logic_vector(23 DOWNTO 0);SIGNAL zed22165f2:std_logic_vector(23 DOWNTO 0);SIGNAL z90a7dbf30:std_logic_vector(23 DOWNTO 0);SIGNAL zf090fac59:std_logic_vector(7 DOWNTO 0);COMPONENT z_black_box_v PORT(clk:IN std_logic ;z28c1a03db:IN std_logic ;zf1caf1a47:IN std_logic_vector(23 DOWNTO 0);rst_n:IN std_logic ;write:IN std_logic ;zaaac8007d:IN std_logic_vector(7 DOWNTO 0);z3417d2827:OUT std_logic_vector(23 DOWNTO 0));END COMPONENT;FOR ALL:z_black_box_v USE ENTITY pre_made.z_black_box_v;BEGIN z508ec0017<=write AND z1934d98a3;zb48298c48<=write AND z0068e7d64;z75dc1577a<=write AND zb30429bb4;z833ab3bd5<=write AND z9f041aaff;zc57c46db4<=write AND zcf058ee7c;z1ea89dc0d<=write AND ze6d31b4ac;zcd48e1f4f<=write AND z1b791bfd5;z36424fa31<=write AND z45a1dff88;z22f92b4dd<='1';zd4351336a:PROCESS(z22f92b4dd, z2677755d9)BEGIN IF(z2677755d9(0)=z22f92b4dd)THEN z36f79a239<="0000";ELSIF(z2677755d9(1)=z22f92b4dd)THEN z36f79a239<="0001";ELSIF(z2677755d9(2)=z22f92b4dd)THEN z36f79a239<="0010";ELSIF(z2677755d9(3)=z22f92b4dd)THEN z36f79a239<="0011";ELSIF(z2677755d9(4)=z22f92b4dd)THEN z36f79a239<="0100";ELSIF(z2677755d9(5)=z22f92b4dd)THEN z36f79a239<="0101";ELSIF(z2677755d9(6)=z22f92b4dd)THEN z36f79a239<="0110";ELSIF(z2677755d9(7)=z22f92b4dd)THEN z36f79a239<="0111";ELSE z36f79a239<="1000";END IF;END PROCESS zd4351336a;zc83e54d35<=z36f79a239(2)& z36f79a239(1)& z36f79a239(0);z16921971f:PROCESS(z3417d2827, z564ee05a3, z0a9315da3, z6bb6c7052, z163c5325c, z84b2eb77e, zed22165f2, z90a7dbf30, zc83e54d35)BEGIN CASE zc83e54d35 IS WHEN"000"=>z921c03197<=z3417d2827;WHEN"001"=>z921c03197<=z564ee05a3;WHEN"010"=>z921c03197<=z0a9315da3;WHEN"011"=>z921c03197<=z6bb6c7052;WHEN"100"=>z921c03197<=z163c5325c;WHEN"101"=>z921c03197<=z84b2eb77e;WHEN"110"=>z921c03197<=zed22165f2;WHEN"111"=>z921c03197<=z90a7dbf30;WHEN OTHERS=>z921c03197<=(OTHERS=>'X');END CASE;END PROCESS z16921971f;zf090fac59<=z2677755d9;z193f2f0f4:PROCESS(zf090fac59)VARIABLE z925f2bf10:std_logic_vector(7 DOWNTO 0);BEGIN z925f2bf10:=zf090fac59(7 DOWNTO 0);z1934d98a3<=z925f2bf10(0);z0068e7d64<=z925f2bf10(1);zb30429bb4<=z925f2bf10(2);z9f041aaff<=z925f2bf10(3);zcf058ee7c<=z925f2bf10(4);ze6d31b4ac<=z925f2bf10(5);z1b791bfd5<=z925f2bf10(6);z45a1dff88<=z925f2bf10(7);END PROCESS z193f2f0f4;U_0:z_black_box_v PORT MAP(clk=>clk,z28c1a03db=>z28c1a03db,zf1caf1a47=>zd58ce0c39,rst_n=>rst_n,write=>z508ec0017,zaaac8007d=>zaaac8007d,z3417d2827=>z3417d2827);U_1:z_black_box_v PORT MAP(clk=>clk,z28c1a03db=>z28c1a03db,zf1caf1a47=>zd58ce0c39,rst_n=>rst_n,write=>zb48298c48,zaaac8007d=>zaaac8007d,z3417d2827=>z564ee05a3);U_2:z_black_box_v PORT MAP(clk=>clk,z28c1a03db=>z28c1a03db,zf1caf1a47=>zd58ce0c39,rst_n=>rst_n,write=>z75dc1577a,zaaac8007d=>zaaac8007d,z3417d2827=>z0a9315da3);U_3:z_black_box_v PORT MAP(clk=>clk,z28c1a03db=>z28c1a03db,zf1caf1a47=>zd58ce0c39,rst_n=>rst_n,write=>z833ab3bd5,zaaac8007d=>zaaac8007d,z3417d2827=>z6bb6c7052);U_4:z_black_box_v PORT MAP(clk=>clk,z28c1a03db=>z28c1a03db,zf1caf1a47=>zd58ce0c39,rst_n=>rst_n,write=>zc57c46db4,zaaac8007d=>zaaac8007d,z3417d2827=>z163c5325c);U_5:z_black_box_v PORT MAP(clk=>clk,z28c1a03db=>z28c1a03db,zf1caf1a47=>zd58ce0c39,rst_n=>rst_n,write=>z1ea89dc0d,zaaac8007d=>zaaac8007d,z3417d2827=>z84b2eb77e);U_6:z_black_box_v PORT MAP(clk=>clk,z28c1a03db=>z28c1a03db,zf1caf1a47=>zd58ce0c39,rst_n=>rst_n,write=>zcd48e1f4f,zaaac8007d=>zaaac8007d,z3417d2827=>zed22165f2);U_7:z_black_box_v PORT MAP(clk=>clk,z28c1a03db=>z28c1a03db,zf1caf1a47=>zd58ce0c39,rst_n=>rst_n,write=>z36424fa31,zaaac8007d=>zaaac8007d,z3417d2827=>z90a7dbf30);END struct;