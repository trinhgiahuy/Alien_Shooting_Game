--* ><(((('> * Puli puli * ><(((('> // Ƹ̵̡Ӝ̵̨̄Ʒ * swish swish* Ƹ̵̡Ӝ̵̨̄Ʒ Ƹ̵̡Ӝ̵̨̄Ʒ // (っ◕‿◕)╭∩╮^H^H^Hっ
LIBRARY ieee;USE ieee.std_logic_1164.all;USE ieee.std_logic_arith.all;ENTITY z_black_box_j IS PORT(clk:IN std_logic;rst_n:IN std_logic;z1c78dfa64:IN std_logic;zea9c5ae7c:OUT std_logic;zc2cbe183e:OUT std_logic;z7975aa26e:OUT std_logic;z2ebb22097:OUT std_logic);END z_black_box_j ;LIBRARY ieee;USE ieee.std_logic_1164.all;USE ieee.std_logic_arith.all;LIBRARY pre_made;ARCHITECTURE struct OF z_black_box_j IS SIGNAL z6168e6eca:std_logic;SIGNAL z7f53ee971:std_logic;COMPONENT z_black_box_s PORT(clk:IN std_logic ;rst_n:IN std_logic ;z7f53ee971:IN std_logic ;zea9c5ae7c:OUT std_logic ;z7975aa26e:OUT std_logic ;z2ebb22097:OUT std_logic);END COMPONENT;COMPONENT z_black_box_t PORT(clk:IN std_logic ;rst_n:IN std_logic ;z6168e6eca:OUT std_logic ;zc2cbe183e:OUT std_logic);END COMPONENT;FOR ALL:z_black_box_s USE ENTITY pre_made.z_black_box_s;FOR ALL:z_black_box_t USE ENTITY pre_made.z_black_box_t;BEGIN z7f53ee971<=z6168e6eca AND z1c78dfa64;U_1:z_black_box_s PORT MAP(clk=>clk,rst_n=>rst_n,z7f53ee971=>z7f53ee971,zea9c5ae7c=>zea9c5ae7c,z7975aa26e=>z7975aa26e,z2ebb22097=>z2ebb22097);U_0:z_black_box_t PORT MAP(clk=>clk,rst_n=>rst_n,z6168e6eca=>z6168e6eca,zc2cbe183e=>zc2cbe183e);END struct;